module forward_unit(
	input wire [4:0] rs1_ex,
	input wire [4:0] rs2_ex,
	input wire [4:0] rd_mem,
	input wire [4:0] rd_wb,
		
	output wire [1:0] mux_alu_1,
	output wire [1:0] mux_alu_2
);

endmodule
